`timescale 1ns / 1ps

module OLEDText(
    );


endmodule
